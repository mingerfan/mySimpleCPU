`define R_OP 7'b011_0011
`define I_OP 7'b000_0011
`define S_OP 7'd010_0011
`define J_OP 7'd110_1111
`define IMM_OP 7'd001_0011
`define LUI_OP 7'd011_0111


`deifne R_FUN7_ADD 7'b000_0000
`define R_FUN7_SUB 7'b010_0000


`define R_FUN3_ADD 3'b000
`define R_FUN3_SUB 3'b000

`define I_FUN3_LW 3'b010

`define IMM_FUN3_ADDI 3'b000

`define S_FUN3_SW 3'd010